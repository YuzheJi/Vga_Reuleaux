module tb_syn_reuleaux();


endmodule: tb_syn_reuleaux
